template_map_withbram.vhd